module sigmoid(
	input [16:0] in,
	output reg [16:0] out
);

integer total;

always @ (in) begin
	case (in)
		17'b01111111111111111: out <= 17'b01111111111111111; //16
		17'b00111111111111111: out <= 17'b01111111111111111; //15
		17'b00011111111111111: out <= 17'b01111111111111111; //14
		17'b00001111111111111: out <= 17'b01111111111111111; //13
		17'b00000111111111111: out <= 17'b01111111111111111; //12
		17'b00000011111111111: out <= 17'b01111111111111111; //11
		17'b00000001111111111: out <= 17'b01111111111111111; //10
		17'b00000000111111111: out <= 17'b01111111111111111; //9
		17'b00000000011111111: out <= 17'b01111111111111111; //8
		17'b00000000001111111: out <= 17'b01111111111111111; //7
		17'b00000000000111111: out <= 17'b01111111111111111; //6
		17'b00000000000011111: out <= 17'b01111111111111111; //5
		17'b00000000000001111: out <= 17'b01111111111111111; //4
		17'b00000000000000111: out <= 17'b00111111111111111; //3
		17'b00000000000000011: out <= 17'b00011111111111111; //2
		17'b00000000000000001: out <= 17'b00000111111111111; //1
		17'b00000000000000000: out <= 17'b00000000011111111; //0
		17'b10000000000000001: out <= 17'b00000000000001111; //-1
		17'b10000000000000011: out <= 17'b00000000000000011; //-2
		17'b10000000000000111: out <= 17'b00000000000000001; //-3
		17'b10000000000001111: out <= 17'b00000000000000000; //-4
		17'b10000000000011111: out <= 17'b00000000000000000; //-5
		17'b10000000000111111: out <= 17'b00000000000000000; //-6
		17'b10000000001111111: out <= 17'b00000000000000000; //-7
		17'b10000000011111111: out <= 17'b00000000000000000; //-8
		17'b10000000111111111: out <= 17'b00000000000000000; //-9
		17'b10000001111111111: out <= 17'b00000000000000000; //-10
		17'b10000011111111111: out <= 17'b00000000000000000; //-11
		17'b10000111111111111: out <= 17'b00000000000000000; //-12
		17'b10001111111111111: out <= 17'b00000000000000000; //-13
		17'b10011111111111111: out <= 17'b00000000000000000; //-14
		17'b10111111111111111: out <= 17'b00000000000000000; //-15
		17'b11111111111111111: out <= 17'b00000000000000000; //-16
	endcase
end

endmodule